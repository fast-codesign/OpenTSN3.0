////////////////////////////////////////////////////////////////////////////
// Verilog module name - sgmii_eth_substitute.v
// Version: SES_V1.0
///////////////////////////////////////////////////////////////////////////
// Description:
//         the file to substitute of sgmii IP core 
///////////////////////////////////////////////////////////////////////////

`timescale 1 ps / 1 ps
module sgmii_eth_substitute (
		input  wire        clk,            
		input  wire        reset,          
		input  wire        ref_clk,        
        
		input  wire        rxp_0,            
		output wire        txp_0,            
		input  wire [4:0]  reg_addr_0,       
		output wire [15:0] reg_data_out_0,   
		input  wire        reg_rd_0,         
		input  wire [15:0] reg_data_in_0,    
		input  wire        reg_wr_0,         
		output wire        reg_busy_0,       
		output wire        tx_clk_0,         
		output wire        rx_clk_0,         
		input  wire        reset_tx_clk_0,   
		input  wire        reset_rx_clk_0,   
		output wire        gmii_rx_dv_0,     
		output wire [7:0]  gmii_rx_d_0,      
		output wire        gmii_rx_err_0,    
		input  wire        gmii_tx_en_0,     
		input  wire [7:0]  gmii_tx_d_0,      
		input  wire        gmii_tx_err_0,    
		output wire        led_crs_0,        
		output wire        led_link_0,       
		output wire        led_panel_link_0, 
		output wire        led_col_0,        
		output wire        led_an_0,         
		output wire        led_char_err_0,   
		output wire        led_disp_err_0,   
		output wire        rx_recovclkout_0, 
        
        input  wire        rxp_1,            
		output wire        txp_1,            
		input  wire [4:0]  reg_addr_1,       
		output wire [15:0] reg_data_out_1,   
		input  wire        reg_rd_1,         
		input  wire [15:0] reg_data_in_1,    
		input  wire        reg_wr_1,         
		output wire        reg_busy_1,       
		output wire        tx_clk_1,         
		output wire        rx_clk_1,         
		input  wire        reset_tx_clk_1,   
		input  wire        reset_rx_clk_1,   
		output wire        gmii_rx_dv_1,     
		output wire [7:0]  gmii_rx_d_1,      
		output wire        gmii_rx_err_1,    
		input  wire        gmii_tx_en_1,     
		input  wire [7:0]  gmii_tx_d_1,      
		input  wire        gmii_tx_err_1,    
		output wire        led_crs_1,        
		output wire        led_link_1,       
		output wire        led_panel_link_1, 
		output wire        led_col_1,        
		output wire        led_an_1,         
		output wire        led_char_err_1,   
		output wire        led_disp_err_1,   
		output wire        rx_recovclkout_1, 
        
        input  wire        rxp_2,            
		output wire        txp_2,            
		input  wire [4:0]  reg_addr_2,       
		output wire [15:0] reg_data_out_2,   
		input  wire        reg_rd_2,         
		input  wire [15:0] reg_data_in_2,    
		input  wire        reg_wr_2,         
		output wire        reg_busy_2,       
		output wire        tx_clk_2,         
		output wire        rx_clk_2,         
		input  wire        reset_tx_clk_2,   
		input  wire        reset_rx_clk_2,   
		output wire        gmii_rx_dv_2,     
		output wire [7:0]  gmii_rx_d_2,      
		output wire        gmii_rx_err_2,    
		input  wire        gmii_tx_en_2,     
		input  wire [7:0]  gmii_tx_d_2,      
		input  wire        gmii_tx_err_2,    
		output wire        led_crs_2,        
		output wire        led_link_2,       
		output wire        led_panel_link_2, 
		output wire        led_col_2,        
		output wire        led_an_2,         
		output wire        led_char_err_2,   
		output wire        led_disp_err_2,   
		output wire        rx_recovclkout_2, 
        
		input  wire        rxp_3,            
		output wire        txp_3,            
		input  wire [4:0]  reg_addr_3,       
		output wire [15:0] reg_data_out_3,   
		input  wire        reg_rd_3,         
		input  wire [15:0] reg_data_in_3,    
		input  wire        reg_wr_3,         
		output wire        reg_busy_3,       
		output wire        tx_clk_3,         
		output wire        rx_clk_3,         
		input  wire        reset_tx_clk_3,   
		input  wire        reset_rx_clk_3,   
		output wire        gmii_rx_dv_3,     
		output wire [7:0]  gmii_rx_d_3,      
		output wire        gmii_rx_err_3,    
		input  wire        gmii_tx_en_3,     
		input  wire [7:0]  gmii_tx_d_3,      
		input  wire        gmii_tx_err_3,    
		output wire        led_crs_3,        
		output wire        led_link_3,       
		output wire        led_panel_link_3, 
		output wire        led_col_3,        
		output wire        led_an_3,         
		output wire        led_char_err_3,   
		output wire        led_disp_err_3,   
		output wire        rx_recovclkout_3  
	);

	wire         i_lvdsio_terminator_0_lvds_rx_inclock_export;                         
	wire  [39:0] i_lvdsio_rx_0_rx_out_export;                                          
	wire   [3:0] i_lvdsio_terminator_0_rx_in_export;                                   
	wire   [3:0] i_lvdsio_terminator_0_rx_dpa_reset_export;                            
	wire   [3:0] i_lvdsio_rx_0_rx_dpa_locked_export;                                   
	wire   [3:0] i_lvdsio_rx_0_rx_divfwdclk_export;                                    
	wire         i_lvdsio_rx_0_rx_coreclock_export;                                    
	wire         i_lvdsio_rx_0_pll_locked_export;                                      
	wire         i_lvdsio_terminator_0_pll_areset_rx_export;                           
	wire         i_lvdsio_terminator_0_lvds_tx_inclock_export;                         
	wire  [39:0] i_lvdsio_terminator_0_tx_in_export;                                   
	wire   [3:0] i_lvdsio_tx_0_tx_out_export;                                          
	wire         i_lvdsio_tx_0_pll_locked_export;                                      
	wire         i_lvdsio_terminator_0_pll_areset_tx_export; 
    
	wire  [9:0] i_tse_pcs_0_tbi_tx_d_muxed_tbi_tx_d_muxed;                             
	wire  [9:0] i_lvdsio_terminator_0_tbi_rx_d_lvds_0_tbi_rx_d_lvds;                   
	wire        i_lvdsio_terminator_0_tbi_rx_clk_0_tbi_rx_clk;                         
	wire        i_lvdsio_terminator_0_rx_reset_sequence_done_0_rx_reset_sequence_done; 
	wire        i_lvdsio_terminator_0_rx_reset_0_rx_reset;                             
	wire        i_lvdsio_terminator_0_tx_reset_0_tx_reset;                             
    
	wire  [9:0] i_tse_pcs_1_tbi_tx_d_muxed_tbi_tx_d_muxed;                             
	wire  [9:0] i_lvdsio_terminator_0_tbi_rx_d_lvds_1_tbi_rx_d_lvds;                   
	wire        i_lvdsio_terminator_0_tbi_rx_clk_1_tbi_rx_clk;                         
	wire        i_lvdsio_terminator_0_rx_reset_sequence_done_1_rx_reset_sequence_done; 
	wire        i_lvdsio_terminator_0_rx_reset_1_rx_reset;                             
	wire        i_lvdsio_terminator_0_tx_reset_1_tx_reset;                             
    
	wire  [9:0] i_tse_pcs_2_tbi_tx_d_muxed_tbi_tx_d_muxed;                             
	wire  [9:0] i_lvdsio_terminator_0_tbi_rx_d_lvds_2_tbi_rx_d_lvds;                   
	wire        i_lvdsio_terminator_0_tbi_rx_clk_2_tbi_rx_clk;                         
	wire        i_lvdsio_terminator_0_rx_reset_sequence_done_2_rx_reset_sequence_done; 
	wire        i_lvdsio_terminator_0_rx_reset_2_rx_reset;                             
	wire        i_lvdsio_terminator_0_tx_reset_2_tx_reset;                             
    
	wire  [9:0] i_tse_pcs_3_tbi_tx_d_muxed_tbi_tx_d_muxed;                             
	wire  [9:0] i_lvdsio_terminator_0_tbi_rx_d_lvds_3_tbi_rx_d_lvds;                   
	wire        i_lvdsio_terminator_0_tbi_rx_clk_3_tbi_rx_clk;                         
	wire        i_lvdsio_terminator_0_rx_reset_sequence_done_3_rx_reset_sequence_done; 
	wire        i_lvdsio_terminator_0_rx_reset_3_rx_reset;                             
	wire        i_lvdsio_terminator_0_tx_reset_3_tx_reset;                             
    
	wire        rst_controller_reset_out_reset;                                        

	altera_eth_tse_pcs_pma_nf_lvds #(
		.ENABLE_TIMESTAMPING (0),
		.DEV_VERSION         (4865),
		.ENABLE_ECC          (0),
		.ENABLE_REV_LOOPBACK (0),
		.DEVICE_FAMILY       ("ARRIA10"),
		.SYNCHRONIZER_DEPTH  (3),
		.ENABLE_CLK_SHARING  (1),
		.ENABLE_SGMII        (0),
		.PHY_IDENTIFIER      (0)
	) i_tse_pcs_0 (
		.clk                    (clk),                                                                  
		.reset                  (reset),                                                                
		.reg_addr               (reg_addr_0),                                                           
		.reg_data_out           (reg_data_out_0),                                                       
		.reg_rd                 (reg_rd_0),                                                             
		.reg_data_in            (reg_data_in_0),                                                        
		.reg_wr                 (reg_wr_0),                                                             
		.reg_busy               (reg_busy_0),                                                           
		.ref_clk                (ref_clk),                                                              
		.gmii_rx_dv             (gmii_rx_dv_0),                                                         
		.gmii_rx_d              (gmii_rx_d_0),                                                          
		.gmii_rx_err            (gmii_rx_err_0),                                                        
		.gmii_tx_en             (gmii_tx_en_0),                                                         
		.gmii_tx_d              (gmii_tx_d_0),                                                          
		.gmii_tx_err            (gmii_tx_err_0),                                                        
		.tx_clk                 (tx_clk_0),                                                             
		.rx_clk                 (rx_clk_0),                                                             
		.reset_tx_clk           (reset_tx_clk_0),                                                       
		.reset_rx_clk           (reset_rx_clk_0),                                                       
		.led_crs                (led_crs_0),                                                            
		.led_link               (led_link_0),                                                           
		.led_panel_link         (led_panel_link_0),                                                     
		.led_col                (led_col_0),                                                            
		.led_an                 (led_an_0),                                                             
		.led_char_err           (led_char_err_0),                                                       
		.led_disp_err           (led_disp_err_0),                                                       
		.rx_recovclkout         (rx_recovclkout_0),                                                     
        
		.rx_reset               (i_lvdsio_terminator_0_rx_reset_0_rx_reset),                            
		.rx_reset_sequence_done (i_lvdsio_terminator_0_rx_reset_sequence_done_0_rx_reset_sequence_done),
		.tbi_rx_clk             (i_lvdsio_terminator_0_tbi_rx_clk_0_tbi_rx_clk),                        
		.tx_reset               (i_lvdsio_terminator_0_tx_reset_0_tx_reset),                            
		.tbi_tx_d_muxed         (i_tse_pcs_0_tbi_tx_d_muxed_tbi_tx_d_muxed),                            
		.tbi_rx_d_lvds          (i_lvdsio_terminator_0_tbi_rx_d_lvds_0_tbi_rx_d_lvds),                  
        
		.tx_clkena              (),                                                                     
		.rx_clkena              (),                                                                     
		.mii_rx_dv              (),                                                                     
		.mii_rx_d               (),                                                                     
		.mii_rx_err             (),                                                                     
		.mii_tx_en              (1'b0),                                                                 
		.mii_tx_d               (4'b0000),                                                              
		.mii_tx_err             (1'b0),                                                                 
		.mii_col                (),                                                                     
		.mii_crs                (),                                                                     
		.set_10                 (),                                                                     
		.set_1000               (),                                                                     
		.set_100                (),                                                                     
		.hd_ena                 (),                                                                     
		.pcs_phase_measure_clk  (1'b0),                                                                 
		.rx_latency_adj         (),                                                                     
		.tx_latency_adj         (),                                                                     
		.tx_ptp_alignment       (),                                                                     
		.pcs_eccstatus          ()                                                                      
	);

	altera_eth_tse_pcs_pma_nf_lvds #(
		.ENABLE_TIMESTAMPING (0),
		.DEV_VERSION         (4865),
		.ENABLE_ECC          (0),
		.ENABLE_REV_LOOPBACK (0),
		.DEVICE_FAMILY       ("ARRIA10"),
		.SYNCHRONIZER_DEPTH  (3),
		.ENABLE_CLK_SHARING  (1),
		.ENABLE_SGMII        (0),
		.PHY_IDENTIFIER      (0)
	) i_tse_pcs_1 (
		.clk                    (clk),                                                                  
		.reset                  (reset),                                                                
		.reg_addr               (reg_addr_1),                                                           
		.reg_data_out           (reg_data_out_1),                                                       
		.reg_rd                 (reg_rd_1),                                                             
		.reg_data_in            (reg_data_in_1),                                                        
		.reg_wr                 (reg_wr_1),                                                             
		.reg_busy               (reg_busy_1),                                                           
		.ref_clk                (ref_clk),                                                              
		.gmii_rx_dv             (gmii_rx_dv_1),                                                         
		.gmii_rx_d              (gmii_rx_d_1),                                                          
		.gmii_rx_err            (gmii_rx_err_1),                                                        
		.gmii_tx_en             (gmii_tx_en_1),                                                         
		.gmii_tx_d              (gmii_tx_d_1),                                                          
		.gmii_tx_err            (gmii_tx_err_1),                                                        
		.tx_clk                 (tx_clk_1),                                                             
		.rx_clk                 (rx_clk_1),                                                             
		.reset_tx_clk           (reset_tx_clk_1),                                                       
		.reset_rx_clk           (reset_rx_clk_1),                                                       
		.led_crs                (led_crs_1),                                                            
		.led_link               (led_link_1),                                                           
		.led_panel_link         (led_panel_link_1),                                                     
		.led_col                (led_col_1),                                                            
		.led_an                 (led_an_1),                                                             
		.led_char_err           (led_char_err_1),                                                       
		.led_disp_err           (led_disp_err_1),                                                       
		.rx_recovclkout         (rx_recovclkout_1),                                                     
        
		.rx_reset               (i_lvdsio_terminator_0_rx_reset_1_rx_reset),                            
		.rx_reset_sequence_done (i_lvdsio_terminator_0_rx_reset_sequence_done_1_rx_reset_sequence_done),
		.tbi_rx_clk             (i_lvdsio_terminator_0_tbi_rx_clk_1_tbi_rx_clk),                        
		.tx_reset               (i_lvdsio_terminator_0_tx_reset_1_tx_reset),                            
		.tbi_tx_d_muxed         (i_tse_pcs_1_tbi_tx_d_muxed_tbi_tx_d_muxed),                            
		.tbi_rx_d_lvds          (i_lvdsio_terminator_0_tbi_rx_d_lvds_1_tbi_rx_d_lvds),                  
        
		.tx_clkena              (),                                                                     
		.rx_clkena              (),                                                                     
		.mii_rx_dv              (),                                                                     
		.mii_rx_d               (),                                                                     
		.mii_rx_err             (),                                                                     
		.mii_tx_en              (1'b0),                                                                 
		.mii_tx_d               (4'b0000),                                                              
		.mii_tx_err             (1'b0),                                                                 
		.mii_col                (),                                                                     
		.mii_crs                (),                                                                     
		.set_10                 (),                                                                     
		.set_1000               (),                                                                     
		.set_100                (),                                                                     
		.hd_ena                 (),                                                                     
		.pcs_phase_measure_clk  (1'b0),                                                                 
		.rx_latency_adj         (),                                                                     
		.tx_latency_adj         (),                                                                     
		.tx_ptp_alignment       (),                                                                     
		.pcs_eccstatus          ()                                                                      
	);
    
    altera_eth_tse_pcs_pma_nf_lvds #(
		.ENABLE_TIMESTAMPING (0),
		.DEV_VERSION         (4865),
		.ENABLE_ECC          (0),
		.ENABLE_REV_LOOPBACK (0),
		.DEVICE_FAMILY       ("ARRIA10"),
		.SYNCHRONIZER_DEPTH  (3),
		.ENABLE_CLK_SHARING  (1),
		.ENABLE_SGMII        (0),
		.PHY_IDENTIFIER      (0)
	) i_tse_pcs_2 (
		.clk                    (clk),                                                                  
		.reset                  (reset),                                                                
		.reg_addr               (reg_addr_2),                                                           
		.reg_data_out           (reg_data_out_2),                                                       
		.reg_rd                 (reg_rd_2),                                                             
		.reg_data_in            (reg_data_in_2),                                                        
		.reg_wr                 (reg_wr_2),                                                             
		.reg_busy               (reg_busy_2),                                                           
		.ref_clk                (ref_clk),                                                              
		.gmii_rx_dv             (gmii_rx_dv_2),                                                         
		.gmii_rx_d              (gmii_rx_d_2),                                                          
		.gmii_rx_err            (gmii_rx_err_2),                                                        
		.gmii_tx_en             (gmii_tx_en_2),                                                         
		.gmii_tx_d              (gmii_tx_d_2),                                                          
		.gmii_tx_err            (gmii_tx_err_2),                                                        
		.tx_clk                 (tx_clk_2),                                                             
		.rx_clk                 (rx_clk_2),                                                             
		.reset_tx_clk           (reset_tx_clk_2),                                                       
		.reset_rx_clk           (reset_rx_clk_2),                                                       
		.led_crs                (led_crs_2),                                                            
		.led_link               (led_link_2),                                                           
		.led_panel_link         (led_panel_link_2),                                                     
		.led_col                (led_col_2),                                                            
		.led_an                 (led_an_2),                                                             
		.led_char_err           (led_char_err_2),                                                       
		.led_disp_err           (led_disp_err_2),                                                       
		.rx_recovclkout         (rx_recovclkout_2),                                                     
        
		.rx_reset               (i_lvdsio_terminator_0_rx_reset_2_rx_reset),                            
		.rx_reset_sequence_done (i_lvdsio_terminator_0_rx_reset_sequence_done_2_rx_reset_sequence_done),
		.tbi_rx_clk             (i_lvdsio_terminator_0_tbi_rx_clk_2_tbi_rx_clk),                        
		.tx_reset               (i_lvdsio_terminator_0_tx_reset_2_tx_reset),                            
		.tbi_tx_d_muxed         (i_tse_pcs_2_tbi_tx_d_muxed_tbi_tx_d_muxed),                            
		.tbi_rx_d_lvds          (i_lvdsio_terminator_0_tbi_rx_d_lvds_2_tbi_rx_d_lvds),                  
        
		.tx_clkena              (),                                                                     
		.rx_clkena              (),                                                                     
		.mii_rx_dv              (),                                                                     
		.mii_rx_d               (),                                                                     
		.mii_rx_err             (),                                                                     
		.mii_tx_en              (1'b0),                                                                 
		.mii_tx_d               (4'b0000),                                                              
		.mii_tx_err             (1'b0),                                                                 
		.mii_col                (),                                                                     
		.mii_crs                (),                                                                     
		.set_20                 (),                                                                     
		.set_2000               (),                                                                     
		.set_200                (),                                                                     
		.hd_ena                 (),                                                                     
		.pcs_phase_measure_clk  (1'b0),                                                                 
		.rx_latency_adj         (),                                                                     
		.tx_latency_adj         (),                                                                     
		.tx_ptp_alignment       (),                                                                     
		.pcs_eccstatus          ()                                                                      
	);

	altera_eth_tse_pcs_pma_nf_lvds #(
		.ENABLE_TIMESTAMPING (0),
		.DEV_VERSION         (4865),
		.ENABLE_ECC          (0),
		.ENABLE_REV_LOOPBACK (0),
		.DEVICE_FAMILY       ("ARRIA10"),
		.SYNCHRONIZER_DEPTH  (3),
		.ENABLE_CLK_SHARING  (1),
		.ENABLE_SGMII        (0),
		.PHY_IDENTIFIER      (0)
	) i_tse_pcs_3 (
		.clk                    (clk),                                                                   
		.reset                  (reset),                                                                 
		.reg_addr               (reg_addr_3),                                                            
		.reg_data_out           (reg_data_out_3),                                                        
		.reg_rd                 (reg_rd_3),                                                              
		.reg_data_in            (reg_data_in_3),                                                         
		.reg_wr                 (reg_wr_3),                                                              
		.reg_busy               (reg_busy_3),                                                            
		.ref_clk                (ref_clk),                                                               
		.gmii_rx_dv             (gmii_rx_dv_3),                                                          
		.gmii_rx_d              (gmii_rx_d_3),                                                           
		.gmii_rx_err            (gmii_rx_err_3),                                                         
		.gmii_tx_en             (gmii_tx_en_3),                                                          
		.gmii_tx_d              (gmii_tx_d_3),                                                           
		.gmii_tx_err            (gmii_tx_err_3),                                                         
		.tx_clk                 (tx_clk_3),                                                              
		.rx_clk                 (rx_clk_3),                                                              
		.reset_tx_clk           (reset_tx_clk_3),                                                        
		.reset_rx_clk           (reset_rx_clk_3),                                                        
		.led_crs                (led_crs_3),                                                             
		.led_link               (led_link_3),                                                            
		.led_panel_link         (led_panel_link_3),                                                      
		.led_col                (led_col_3),                                                             
		.led_an                 (led_an_3),                                                              
		.led_char_err           (led_char_err_3),                                                        
		.led_disp_err           (led_disp_err_3),                                                        
		.rx_recovclkout         (rx_recovclkout_3),                                                      
        
		.rx_reset               (i_lvdsio_terminator_0_rx_reset_3_rx_reset),                             
		.rx_reset_sequence_done (i_lvdsio_terminator_0_rx_reset_sequence_done_3_rx_reset_sequence_done), 
		.tbi_rx_clk             (i_lvdsio_terminator_0_tbi_rx_clk_3_tbi_rx_clk),                         
		.tx_reset               (i_lvdsio_terminator_0_tx_reset_3_tx_reset),                             
		.tbi_tx_d_muxed         (i_tse_pcs_3_tbi_tx_d_muxed_tbi_tx_d_muxed),                             
		.tbi_rx_d_lvds          (i_lvdsio_terminator_0_tbi_rx_d_lvds_3_tbi_rx_d_lvds),                   
        
		.tx_clkena              (),                                                                      
		.rx_clkena              (),                                                                      
		.mii_rx_dv              (),                                                                      
		.mii_rx_d               (),                                                                      
		.mii_rx_err             (),                                                                      
		.mii_tx_en              (1'b0),                                                                  
		.mii_tx_d               (4'b0000),                                                               
		.mii_tx_err             (1'b0),                                                                  
		.mii_col                (),                                                                      
		.mii_crs                (),                                                                      
		.set_30                 (),                                                                      
		.set_3000               (),                                                                      
		.set_300                (),                                                                      
		.hd_ena                 (),                                                                      
		.pcs_phase_measure_clk  (1'b0),                                                                  
		.rx_latency_adj         (),                                                                      
		.tx_latency_adj         (),                                                                      
		.tx_ptp_alignment       (),                                                                      
		.pcs_eccstatus          ()                                                                       
	);
    
	sgmii_pcs_share_altera_lvds_191_xvdv7pi i_lvdsio_rx_0 (
		.rx_in         (i_lvdsio_terminator_0_rx_in_export),          
		.rx_out        (i_lvdsio_rx_0_rx_out_export),                 
		.rx_coreclock  (i_lvdsio_rx_0_rx_coreclock_export),           
		.inclock       (i_lvdsio_terminator_0_lvds_rx_inclock_export),
		.pll_areset    (i_lvdsio_terminator_0_pll_areset_rx_export),  
		.rx_dpa_locked (i_lvdsio_rx_0_rx_dpa_locked_export),          
		.rx_dpa_reset  (i_lvdsio_terminator_0_rx_dpa_reset_export),   
		.rx_divfwdclk  (i_lvdsio_rx_0_rx_divfwdclk_export),           
		.pll_locked    (i_lvdsio_rx_0_pll_locked_export)              
	);

	sgmii_pcs_share_altera_lvds_191_id6gcay i_lvdsio_tx_0 (
		.tx_in      (i_lvdsio_terminator_0_tx_in_export),           
		.tx_out     (i_lvdsio_tx_0_tx_out_export),                  
		.inclock    (i_lvdsio_terminator_0_lvds_tx_inclock_export), 
		.pll_areset (i_lvdsio_terminator_0_pll_areset_tx_export),   
		.pll_locked (i_lvdsio_tx_0_pll_locked_export)               
	);

	altera_eth_tse_nf_lvds_terminator #(
		.NUM_CHANNELS       (4),
		.SYNCHRONIZER_DEPTH (3)
	) i_lvdsio_terminator_0 (
		.lvds_inclock              (ref_clk),                                                              
		.reset                     (rst_controller_reset_out_reset),                                       
		.lvds_rx_inclock           (i_lvdsio_terminator_0_lvds_rx_inclock_export),                         
		.pll_areset_rx             (i_lvdsio_terminator_0_pll_areset_rx_export),                           
		.pll_locked_tx             (i_lvdsio_tx_0_pll_locked_export),                                      
		.lvds_tx_inclock           (i_lvdsio_terminator_0_lvds_tx_inclock_export),                         
		.rx_coreclock              (i_lvdsio_rx_0_rx_coreclock_export),                                    
		.pll_areset_tx             (i_lvdsio_terminator_0_pll_areset_tx_export),                           
		.pll_locked_rx             (i_lvdsio_rx_0_pll_locked_export),                                      
		.rx_dpa_reset              (i_lvdsio_terminator_0_rx_dpa_reset_export),                            
		.rx_in                     (i_lvdsio_terminator_0_rx_in_export),                                   
		.rx_out                    (i_lvdsio_rx_0_rx_out_export),                                          
		.tx_in                     (i_lvdsio_terminator_0_tx_in_export),                                   
		.rx_dpa_locked             (i_lvdsio_rx_0_rx_dpa_locked_export),                                   
		.rx_divfwdclk              (i_lvdsio_rx_0_rx_divfwdclk_export),                                    
		.tx_out                    (i_lvdsio_tx_0_tx_out_export),                                          
        
		.rxp_0                     (rxp_0), 
		.txp_0                     (txp_0), 
		.rx_reset_0                (i_lvdsio_terminator_0_rx_reset_0_rx_reset),                            
		.rx_reset_sequence_done_0  (i_lvdsio_terminator_0_rx_reset_sequence_done_0_rx_reset_sequence_done),
		.tbi_rx_clk_0              (i_lvdsio_terminator_0_tbi_rx_clk_0_tbi_rx_clk),                        
		.tx_reset_0                (i_lvdsio_terminator_0_tx_reset_0_tx_reset),                            
		.tbi_rx_d_lvds_0           (i_lvdsio_terminator_0_tbi_rx_d_lvds_0_tbi_rx_d_lvds),                  
		.tbi_tx_d_muxed_0          (i_tse_pcs_0_tbi_tx_d_muxed_tbi_tx_d_muxed),                            
        
		.rxp_1                     (rxp_1), 
		.txp_1                     (txp_1), 
		.rx_reset_1                (i_lvdsio_terminator_0_rx_reset_1_rx_reset),                            
		.rx_reset_sequence_done_1  (i_lvdsio_terminator_0_rx_reset_sequence_done_1_rx_reset_sequence_done),
		.tbi_rx_clk_1              (i_lvdsio_terminator_0_tbi_rx_clk_1_tbi_rx_clk),                        
		.tx_reset_1                (i_lvdsio_terminator_0_tx_reset_1_tx_reset),                            
		.tbi_rx_d_lvds_1           (i_lvdsio_terminator_0_tbi_rx_d_lvds_1_tbi_rx_d_lvds),                  
		.tbi_tx_d_muxed_1          (i_tse_pcs_1_tbi_tx_d_muxed_tbi_tx_d_muxed),                            
        
		.rxp_2                     (rxp_2), 
		.txp_2                     (txp_2), 
		.rx_reset_2                (i_lvdsio_terminator_0_rx_reset_2_rx_reset),                            
		.rx_reset_sequence_done_2  (i_lvdsio_terminator_0_rx_reset_sequence_done_2_rx_reset_sequence_done),
		.tbi_rx_clk_2              (i_lvdsio_terminator_0_tbi_rx_clk_2_tbi_rx_clk),                        
		.tx_reset_2                (i_lvdsio_terminator_0_tx_reset_2_tx_reset),                            
		.tbi_rx_d_lvds_2           (i_lvdsio_terminator_0_tbi_rx_d_lvds_2_tbi_rx_d_lvds),                  
		.tbi_tx_d_muxed_2          (i_tse_pcs_2_tbi_tx_d_muxed_tbi_tx_d_muxed),                            
        
		.rxp_3                     (rxp_3), 
		.txp_3                     (txp_3), 
		.rx_reset_3                (i_lvdsio_terminator_0_rx_reset_3_rx_reset),                            
		.rx_reset_sequence_done_3  (i_lvdsio_terminator_0_rx_reset_sequence_done_3_rx_reset_sequence_done),
		.tbi_rx_clk_3              (i_lvdsio_terminator_0_tbi_rx_clk_3_tbi_rx_clk),                        
		.tx_reset_3                (i_lvdsio_terminator_0_tx_reset_3_tx_reset),                            
		.tbi_rx_d_lvds_3           (i_lvdsio_terminator_0_tbi_rx_d_lvds_3_tbi_rx_d_lvds),                  
		.tbi_tx_d_muxed_3          (i_tse_pcs_3_tbi_tx_d_muxed_tbi_tx_d_muxed),                            
        
		.rxp_4                     (1'b0),                                                                 
		.txp_4                     (),                                                                     
		.rx_reset_4                (),                                                                     
		.rx_reset_sequence_done_4  (),                                                                     
		.tbi_rx_clk_4              (),                                                                     
		.tx_reset_4                (),                                                                     
		.tbi_rx_d_lvds_4           (),                                                                     
		.tbi_tx_d_muxed_4          (10'b0000000000),                                                       
        
		.rxp_5                     (1'b0),                                                                 
		.txp_5                     (),                                                                     
		.rx_reset_5                (),                                                                     
		.rx_reset_sequence_done_5  (),                                                                     
		.tbi_rx_clk_5              (),                                                                     
		.tx_reset_5                (),                                                                     
		.tbi_rx_d_lvds_5           (),                                                                     
		.tbi_tx_d_muxed_5          (10'b0000000000),                                                       
        
		.rxp_6                     (1'b0),                                                                 
		.txp_6                     (),                                                                     
		.rx_reset_6                (),                                                                     
		.rx_reset_sequence_done_6  (),                                                                     
		.tbi_rx_clk_6              (),                                                                     
		.tx_reset_6                (),                                                                     
		.tbi_rx_d_lvds_6           (),                                                                     
		.tbi_tx_d_muxed_6          (10'b0000000000),                                                       
        
		.rxp_7                     (1'b0),                                                                 
		.txp_7                     (),                                                                     
		.rx_reset_7                (),                                                                     
		.rx_reset_sequence_done_7  (),                                                                     
		.tbi_rx_clk_7              (),                                                                     
		.tx_reset_7                (),                                                                     
		.tbi_rx_d_lvds_7           (),                                                                     
		.tbi_tx_d_muxed_7          (10'b0000000000),                                                       
        
		.rxp_8                     (1'b0),                                                                 
		.txp_8                     (),                                                                     
		.rx_reset_8                (),                                                                     
		.rx_reset_sequence_done_8  (),                                                                     
		.tbi_rx_clk_8              (),                                                                     
		.tx_reset_8                (),                                                                     
		.tbi_rx_d_lvds_8           (),                                                                     
		.tbi_tx_d_muxed_8          (10'b0000000000),                                                       
        
		.rxp_9                     (1'b0),                                                                 
		.txp_9                     (),                                                                     
		.rx_reset_9                (),                                                                     
		.rx_reset_sequence_done_9  (),                                                                     
		.tbi_rx_clk_9              (),                                                                     
		.tx_reset_9                (),                                                                     
		.tbi_rx_d_lvds_9           (),                                                                     
		.tbi_tx_d_muxed_9          (10'b0000000000),                                                       
        
		.rxp_10                    (1'b0),                                                                 
		.txp_10                    (),                                                                     
		.rx_reset_10               (),                                                                     
		.rx_reset_sequence_done_10 (),                                                                     
		.tbi_rx_clk_10             (),                                                                     
		.tx_reset_10               (),                                                                     
		.tbi_rx_d_lvds_10          (),                                                                     
		.tbi_tx_d_muxed_10         (10'b0000000000),                                                       
        
		.rxp_11                    (1'b0),                                                                 
		.txp_11                    (),                                                                     
		.rx_reset_11               (),                                                                     
		.rx_reset_sequence_done_11 (),                                                                     
		.tbi_rx_clk_11             (),                                                                     
		.tx_reset_11               (),                                                                     
		.tbi_rx_d_lvds_11          (),                                                                     
		.tbi_tx_d_muxed_11         (10'b0000000000)                                                        
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (reset),                          
		.clk            (ref_clk),                        
		.reset_out      (rst_controller_reset_out_reset), 
		.reset_req      (),                               
		.reset_req_in0  (1'b0),                           
		.reset_in1      (1'b0),                           
		.reset_req_in1  (1'b0),                           
		.reset_in2      (1'b0),                           
		.reset_req_in2  (1'b0),                           
		.reset_in3      (1'b0),                           
		.reset_req_in3  (1'b0),                           
		.reset_in4      (1'b0),                           
		.reset_req_in4  (1'b0),                           
		.reset_in5      (1'b0),                           
		.reset_req_in5  (1'b0),                           
		.reset_in6      (1'b0),                           
		.reset_req_in6  (1'b0),                           
		.reset_in7      (1'b0),                           
		.reset_req_in7  (1'b0),                           
		.reset_in8      (1'b0),                           
		.reset_req_in8  (1'b0),                           
		.reset_in9      (1'b0),                           
		.reset_req_in9  (1'b0),                           
		.reset_in10     (1'b0),                           
		.reset_req_in10 (1'b0),                           
		.reset_in11     (1'b0),                           
		.reset_req_in11 (1'b0),                           
		.reset_in12     (1'b0),                           
		.reset_req_in12 (1'b0),                           
		.reset_in13     (1'b0),                           
		.reset_req_in13 (1'b0),                           
		.reset_in14     (1'b0),                           
		.reset_req_in14 (1'b0),                           
		.reset_in15     (1'b0),                           
		.reset_req_in15 (1'b0)                            
	);

endmodule
