////////////////////////////////////////////////////////////////////////////
// Verilog module name - sgmii_substitute.v
// Version: SST_V1.0
///////////////////////////////////////////////////////////////////////////
// Description:
//         the file to substitute of sgmii IP core 
///////////////////////////////////////////////////////////////////////////

`timescale 1 ps / 1 ps
module sgmii_substitute (
		input  wire        clk,            
		input  wire        reset,          
		input  wire        ref_clk,        
        
		input  wire        rxp_0,            
		output wire        txp_0,            
		input  wire [4:0]  reg_addr_0,       
		output wire [15:0] reg_data_out_0,   
		input  wire        reg_rd_0,         
		input  wire [15:0] reg_data_in_0,    
		input  wire        reg_wr_0,         
		output wire        reg_busy_0,       
		output wire        tx_clk_0,         
		output wire        rx_clk_0,         
		input  wire        reset_tx_clk_0,   
		input  wire        reset_rx_clk_0,   
		output wire        gmii_rx_dv_0,     
		output wire [7:0]  gmii_rx_d_0,      
		output wire        gmii_rx_err_0,    
		input  wire        gmii_tx_en_0,     
		input  wire [7:0]  gmii_tx_d_0,      
		input  wire        gmii_tx_err_0,    
		output wire        led_crs_0,        
		output wire        led_link_0,       
		output wire        led_panel_link_0, 
		output wire        led_col_0,        
		output wire        led_an_0,         
		output wire        led_char_err_0,   
		output wire        led_disp_err_0,   
		output wire        rx_recovclkout_0, 
        
        input  wire        rxp_1,            
		output wire        txp_1,            
		input  wire [4:0]  reg_addr_1,       
		output wire [15:0] reg_data_out_1,   
		input  wire        reg_rd_1,         
		input  wire [15:0] reg_data_in_1,    
		input  wire        reg_wr_1,         
		output wire        reg_busy_1,       
		output wire        tx_clk_1,         
		output wire        rx_clk_1,         
		input  wire        reset_tx_clk_1,   
		input  wire        reset_rx_clk_1,   
		output wire        gmii_rx_dv_1,    
		output wire [7:0]  gmii_rx_d_1,     
		output wire        gmii_rx_err_1,   
		input  wire        gmii_tx_en_1,    
		input  wire [7:0]  gmii_tx_d_1,     
		input  wire        gmii_tx_err_1,   
		output wire        led_crs_1,       
		output wire        led_link_1,      
		output wire        led_panel_link_1,
		output wire        led_col_1,       
		output wire        led_an_1,        
		output wire        led_char_err_1,  
		output wire        led_disp_err_1,  
		output wire        rx_recovclkout_1,
        
        input  wire        rxp_2,           
		output wire        txp_2,           
		input  wire [4:0]  reg_addr_2,      
		output wire [15:0] reg_data_out_2,  
		input  wire        reg_rd_2,        
		input  wire [15:0] reg_data_in_2,   
		input  wire        reg_wr_2,        
		output wire        reg_busy_2,      
		output wire        tx_clk_2,        
		output wire        rx_clk_2,        
		input  wire        reset_tx_clk_2,  
		input  wire        reset_rx_clk_2,  
		output wire        gmii_rx_dv_2,    
		output wire [7:0]  gmii_rx_d_2,     
		output wire        gmii_rx_err_2,   
		input  wire        gmii_tx_en_2,    
		input  wire [7:0]  gmii_tx_d_2,     
		input  wire        gmii_tx_err_2,   
		output wire        led_crs_2,       
		output wire        led_link_2,      
		output wire        led_panel_link_2,
		output wire        led_col_2,       
		output wire        led_an_2,        
		output wire        led_char_err_2,  
		output wire        led_disp_err_2,  
		output wire        rx_recovclkout_2,
        
		input  wire        rxp_3,           
		output wire        txp_3,           
		input  wire [4:0]  reg_addr_3,      
		output wire [15:0] reg_data_out_3,  
		input  wire        reg_rd_3,        
		input  wire [15:0] reg_data_in_3,   
		input  wire        reg_wr_3,        
		output wire        reg_busy_3,      
		output wire        tx_clk_3,        
		output wire        rx_clk_3,        
		input  wire        reset_tx_clk_3,  
		input  wire        reset_rx_clk_3,  
		output wire        gmii_rx_dv_3,    
		output wire [7:0]  gmii_rx_d_3,     
		output wire        gmii_rx_err_3,   
		input  wire        gmii_tx_en_3,    
		input  wire [7:0]  gmii_tx_d_3,     
		input  wire        gmii_tx_err_3,   
		output wire        led_crs_3,       
		output wire        led_link_3,      
		output wire        led_panel_link_3,
		output wire        led_col_3,       
		output wire        led_an_3,        
		output wire        led_char_err_3,  
		output wire        led_disp_err_3,  
		output wire        rx_recovclkout_3 
	);

	sgmii_eth_substitute eth_tse_0 (
		.clk            (clk),            
		.reset          (reset),          
		.ref_clk        (ref_clk),        
        
		.rxp_0            (rxp_0),            
		.txp_0            (txp_0),            
		.reg_addr_0       (reg_addr_0),       
		.reg_data_out_0   (reg_data_out_0),   
		.reg_rd_0         (reg_rd_0),         
		.reg_data_in_0    (reg_data_in_0),    
		.reg_wr_0         (reg_wr_0),         
		.reg_busy_0       (reg_busy_0),       
		.tx_clk_0         (tx_clk_0),         
		.rx_clk_0         (rx_clk_0),         
		.reset_tx_clk_0   (reset_tx_clk_0),   
		.reset_rx_clk_0   (reset_rx_clk_0),   
		.gmii_rx_dv_0     (gmii_rx_dv_0),     
		.gmii_rx_d_0      (gmii_rx_d_0),      
		.gmii_rx_err_0    (gmii_rx_err_0),    
		.gmii_tx_en_0     (gmii_tx_en_0),     
		.gmii_tx_d_0      (gmii_tx_d_0),      
		.gmii_tx_err_0    (gmii_tx_err_0),    
		.led_crs_0        (led_crs_0),        
		.led_link_0       (led_link_0),       
		.led_panel_link_0 (led_panel_link_0), 
		.led_col_0        (led_col_0),        
		.led_an_0         (led_an_0),         
		.led_char_err_0   (led_char_err_0),   
		.led_disp_err_0   (led_disp_err_0),   
		.rx_recovclkout_0 (rx_recovclkout_0), 
        
		.rxp_1            (rxp_1),            
		.txp_1            (txp_1),            
		.reg_addr_1       (reg_addr_1),       
		.reg_data_out_1   (reg_data_out_1),   
		.reg_rd_1         (reg_rd_1),         
		.reg_data_in_1    (reg_data_in_1),    
		.reg_wr_1         (reg_wr_1),         
		.reg_busy_1       (reg_busy_1),       
		.tx_clk_1         (tx_clk_1),         
		.rx_clk_1         (rx_clk_1),         
		.reset_tx_clk_1   (reset_tx_clk_1),   
		.reset_rx_clk_1   (reset_rx_clk_1),   
		.gmii_rx_dv_1     (gmii_rx_dv_1),     
		.gmii_rx_d_1      (gmii_rx_d_1),      
		.gmii_rx_err_1    (gmii_rx_err_1),    
		.gmii_tx_en_1     (gmii_tx_en_1),     
		.gmii_tx_d_1      (gmii_tx_d_1),      
		.gmii_tx_err_1    (gmii_tx_err_1),    
		.led_crs_1        (led_crs_1),        
		.led_link_1       (led_link_1),       
		.led_panel_link_1 (led_panel_link_1), 
		.led_col_1        (led_col_1),        
		.led_an_1         (led_an_1),         
		.led_char_err_1   (led_char_err_1),   
		.led_disp_err_1   (led_disp_err_1),   
		.rx_recovclkout_1 (rx_recovclkout_1), 
        
        .rxp_2            (rxp_2),            
		.txp_2            (txp_2),            
		.reg_addr_2       (reg_addr_2),       
		.reg_data_out_2   (reg_data_out_2),   
		.reg_rd_2         (reg_rd_2),         
		.reg_data_in_2    (reg_data_in_2),    
		.reg_wr_2         (reg_wr_2),         
		.reg_busy_2       (reg_busy_2),       
		.tx_clk_2         (tx_clk_2),         
		.rx_clk_2         (rx_clk_2),         
		.reset_tx_clk_2   (reset_tx_clk_2),   
		.reset_rx_clk_2   (reset_rx_clk_2),   
		.gmii_rx_dv_2     (gmii_rx_dv_2),     
		.gmii_rx_d_2      (gmii_rx_d_2),      
		.gmii_rx_err_2    (gmii_rx_err_2),    
		.gmii_tx_en_2     (gmii_tx_en_2),     
		.gmii_tx_d_2      (gmii_tx_d_2),      
		.gmii_tx_err_2    (gmii_tx_err_2),    
		.led_crs_2        (led_crs_2),        
		.led_link_2       (led_link_2),       
		.led_panel_link_2 (led_panel_link_2), 
		.led_col_2        (led_col_2),        
		.led_an_2         (led_an_2),         
		.led_char_err_2   (led_char_err_2),   
		.led_disp_err_2   (led_disp_err_2),   
		.rx_recovclkout_2 (rx_recovclkout_2), 
        
        .rxp_3            (rxp_3),            
		.txp_3            (txp_3),            
		.reg_addr_3       (reg_addr_3),       
		.reg_data_out_3   (reg_data_out_3),   
		.reg_rd_3         (reg_rd_3),         
		.reg_data_in_3    (reg_data_in_3),    
		.reg_wr_3         (reg_wr_3),         
		.reg_busy_3       (reg_busy_3),       
		.tx_clk_3         (tx_clk_3),         
		.rx_clk_3         (rx_clk_3),         
		.reset_tx_clk_3   (reset_tx_clk_3),   
		.reset_rx_clk_3   (reset_rx_clk_3),   
		.gmii_rx_dv_3     (gmii_rx_dv_3),     
		.gmii_rx_d_3      (gmii_rx_d_3),      
		.gmii_rx_err_3    (gmii_rx_err_3),    
		.gmii_tx_en_3     (gmii_tx_en_3),     
		.gmii_tx_d_3      (gmii_tx_d_3),      
		.gmii_tx_err_3    (gmii_tx_err_3),    
		.led_crs_3        (led_crs_3),        
		.led_link_3       (led_link_3),       
		.led_panel_link_3 (led_panel_link_3), 
		.led_col_3        (led_col_3),        
		.led_an_3         (led_an_3),         
		.led_char_err_3   (led_char_err_3),   
		.led_disp_err_3   (led_disp_err_3),   
		.rx_recovclkout_3 (rx_recovclkout_3)  
	);

endmodule
